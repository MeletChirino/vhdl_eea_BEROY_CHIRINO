library	ieee;
use	ieee.std_logic_1164.all;
use 	ieee.std_logic_unsigned.all;
use 	ieee.numeric_std.all;

package tools is

	component pwm_module is
		port(
			freq	: in std_logic_vector(15 downto 0);
			duty	: in std_logic_vector(15 downto 0);
			clk_in	: in std_logic;
			pwm	: out std_logic
		    );
	end component;
	component clk_1MHz is
		port(
			clk_in	: in std_logic;
			clk_out	: out std_logic
		    );
	end component;
	component shift_register is
		port(
			data_in		: in std_logic;
			angle_barre	: out std_logic_vector(11 downto 0);
			clk_in		: in std_logic := '0'
		);
	end component;
	component clk_50MHz is
		port(
			output	: out std_logic := 0
	    );
	end component;
end tools;
