-- Filr 
library	ieee;
use	ieee.std_logic_1164.all;
use 	ieee.std_logic_unsigned.all;
use	ieee.numeric_std.all;

--my components
library work;
use	work.tools.all;

entity gestion_verin is
end entity;

architecture rtl of gestion_verin is

begin
	

end rtl;
