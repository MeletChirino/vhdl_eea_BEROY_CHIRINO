
module mon_pwm (
	clk_clk,
	pwm_0_conduit_end_writeresponsevalid_n);	

	input		clk_clk;
	output		pwm_0_conduit_end_writeresponsevalid_n;
endmodule
