  --Example instantiation for system 'MicroAnemo'
  MicroAnemo_inst : MicroAnemo
    port map(
      clk_0 => clk_0,
      in_port_to_the_freq_out => in_port_to_the_freq_out,
      reset_n => reset_n
    );


