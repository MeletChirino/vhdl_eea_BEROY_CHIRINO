-- sopc3.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sopc3 is
	port (
		angle_barre_external_connection_export : out std_logic_vector(11 downto 0);                    -- angle_barre_external_connection.export
		butee_d_external_connection_export     : out std_logic_vector(11 downto 0);                    --     butee_d_external_connection.export
		butee_g_external_connection_export     : out std_logic_vector(11 downto 0);                    --     butee_g_external_connection.export
		clk_clk                                : in  std_logic                     := '0';             --                             clk.clk
		duty_external_connection_export        : out std_logic_vector(15 downto 0);                    --        duty_external_connection.export
		freq_external_connection_export        : out std_logic_vector(15 downto 0);                    --        freq_external_connection.export
		sens_external_connection_export        : out std_logic;                                        --        sens_external_connection.export
		write_data_external_connection_export  : in  std_logic_vector(7 downto 0)  := (others => '0'); --  write_data_external_connection.export
		write_n_external_connection_export     : in  std_logic                     := '0'              --     write_n_external_connection.export
	);
end entity sopc3;

architecture rtl of sopc3 is
	component sopc3_angle_barre is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(11 downto 0)                     -- export
		);
	end component sopc3_angle_barre;

	component sopc3_duty is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component sopc3_duty;

	component sopc3_intel_generic_serial_flash_interface_top_0 is
		generic (
			DEVICE_FAMILY : string  := "";
			CHIP_SELS     : integer := 1
		);
		port (
			avl_csr_address       : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			avl_csr_read          : in  std_logic                     := 'X';             -- read
			avl_csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avl_csr_write         : in  std_logic                     := 'X';             -- write
			avl_csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_csr_waitrequest   : out std_logic;                                        -- waitrequest
			avl_csr_readdatavalid : out std_logic;                                        -- readdatavalid
			avl_mem_write         : in  std_logic                     := 'X';             -- write
			avl_mem_burstcount    : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			avl_mem_waitrequest   : out std_logic;                                        -- waitrequest
			avl_mem_read          : in  std_logic                     := 'X';             -- read
			avl_mem_address       : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			avl_mem_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_mem_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avl_mem_readdatavalid : out std_logic;                                        -- readdatavalid
			avl_mem_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk_clk               : in  std_logic                     := 'X';             -- clk
			reset_reset           : in  std_logic                     := 'X'              -- reset
		);
	end component sopc3_intel_generic_serial_flash_interface_top_0;

	component sopc3_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component sopc3_jtag_uart_0;

	component sopc3_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(23 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(23 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component sopc3_nios2_gen2_0;

	component sopc3_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component sopc3_onchip_memory2_0;

	component sopc3_sens is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component sopc3_sens;

	component sopc3_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component sopc3_sysid_qsys_0;

	component sopc3_write_data is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component sopc3_write_data;

	component sopc3_write_n is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component sopc3_write_n;

	component sopc3_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                                                : in  std_logic                     := 'X';             -- clk
			intel_generic_serial_flash_interface_top_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                               : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                                             : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                                         : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                                                : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                                            : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                                               : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                                         : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                                      : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                                  : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                                         : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                                     : out std_logic_vector(31 downto 0);                    -- readdata
			angle_barre_s1_address                                                       : out std_logic_vector(1 downto 0);                     -- address
			angle_barre_s1_write                                                         : out std_logic;                                        -- write
			angle_barre_s1_readdata                                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			angle_barre_s1_writedata                                                     : out std_logic_vector(31 downto 0);                    -- writedata
			angle_barre_s1_chipselect                                                    : out std_logic;                                        -- chipselect
			butee_d_s1_address                                                           : out std_logic_vector(1 downto 0);                     -- address
			butee_d_s1_write                                                             : out std_logic;                                        -- write
			butee_d_s1_readdata                                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			butee_d_s1_writedata                                                         : out std_logic_vector(31 downto 0);                    -- writedata
			butee_d_s1_chipselect                                                        : out std_logic;                                        -- chipselect
			butee_g_s1_address                                                           : out std_logic_vector(1 downto 0);                     -- address
			butee_g_s1_write                                                             : out std_logic;                                        -- write
			butee_g_s1_readdata                                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			butee_g_s1_writedata                                                         : out std_logic_vector(31 downto 0);                    -- writedata
			butee_g_s1_chipselect                                                        : out std_logic;                                        -- chipselect
			duty_s1_address                                                              : out std_logic_vector(1 downto 0);                     -- address
			duty_s1_write                                                                : out std_logic;                                        -- write
			duty_s1_readdata                                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			duty_s1_writedata                                                            : out std_logic_vector(31 downto 0);                    -- writedata
			duty_s1_chipselect                                                           : out std_logic;                                        -- chipselect
			freq_s1_address                                                              : out std_logic_vector(1 downto 0);                     -- address
			freq_s1_write                                                                : out std_logic;                                        -- write
			freq_s1_readdata                                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			freq_s1_writedata                                                            : out std_logic_vector(31 downto 0);                    -- writedata
			freq_s1_chipselect                                                           : out std_logic;                                        -- chipselect
			intel_generic_serial_flash_interface_top_0_avl_csr_address                   : out std_logic_vector(5 downto 0);                     -- address
			intel_generic_serial_flash_interface_top_0_avl_csr_write                     : out std_logic;                                        -- write
			intel_generic_serial_flash_interface_top_0_avl_csr_read                      : out std_logic;                                        -- read
			intel_generic_serial_flash_interface_top_0_avl_csr_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			intel_generic_serial_flash_interface_top_0_avl_csr_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid             : in  std_logic                     := 'X';             -- readdatavalid
			intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			intel_generic_serial_flash_interface_top_0_avl_mem_address                   : out std_logic_vector(19 downto 0);                    -- address
			intel_generic_serial_flash_interface_top_0_avl_mem_write                     : out std_logic;                                        -- write
			intel_generic_serial_flash_interface_top_0_avl_mem_read                      : out std_logic;                                        -- read
			intel_generic_serial_flash_interface_top_0_avl_mem_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			intel_generic_serial_flash_interface_top_0_avl_mem_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			intel_generic_serial_flash_interface_top_0_avl_mem_burstcount                : out std_logic_vector(6 downto 0);                     -- burstcount
			intel_generic_serial_flash_interface_top_0_avl_mem_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid             : in  std_logic                     := 'X';             -- readdatavalid
			intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_address                                        : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                                          : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                                           : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                                    : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                                     : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                                         : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                                           : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                                            : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                                      : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                                     : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                                     : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                                                  : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s1_write                                                    : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                                               : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                                               : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                                    : out std_logic;                                        -- clken
			sens_s1_address                                                              : out std_logic_vector(1 downto 0);                     -- address
			sens_s1_write                                                                : out std_logic;                                        -- write
			sens_s1_readdata                                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sens_s1_writedata                                                            : out std_logic_vector(31 downto 0);                    -- writedata
			sens_s1_chipselect                                                           : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                                           : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			write_data_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			write_data_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			write_n_s1_address                                                           : out std_logic_vector(1 downto 0);                     -- address
			write_n_s1_readdata                                                          : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component sopc3_mm_interconnect_0;

	component sopc3_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component sopc3_irq_mapper;

	component sopc3_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component sopc3_rst_controller;

	component sopc3_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component sopc3_rst_controller_001;

	signal nios2_gen2_0_debug_reset_request_reset                                             : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_001:reset_in1]
	signal nios2_gen2_0_data_master_readdata                                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                               : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                               : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                                   : std_logic_vector(23 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                                : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                                      : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                                     : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                                 : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                            : std_logic_vector(23 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                               : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect                         : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                           : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest                        : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                               : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                              : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_readdata      : std_logic_vector(31 downto 0); -- intel_generic_serial_flash_interface_top_0:avl_csr_readdata -> mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_csr_readdata
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest   : std_logic;                     -- intel_generic_serial_flash_interface_top_0:avl_csr_waitrequest -> mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_address       : std_logic_vector(5 downto 0);  -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_csr_address -> intel_generic_serial_flash_interface_top_0:avl_csr_address
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_read          : std_logic;                     -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_csr_read -> intel_generic_serial_flash_interface_top_0:avl_csr_read
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid : std_logic;                     -- intel_generic_serial_flash_interface_top_0:avl_csr_readdatavalid -> mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_write         : std_logic;                     -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_csr_write -> intel_generic_serial_flash_interface_top_0:avl_csr_write
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_csr_writedata -> intel_generic_serial_flash_interface_top_0:avl_csr_writedata
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_readdata      : std_logic_vector(31 downto 0); -- intel_generic_serial_flash_interface_top_0:avl_mem_readdata -> mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_mem_readdata
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest   : std_logic;                     -- intel_generic_serial_flash_interface_top_0:avl_mem_waitrequest -> mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_address       : std_logic_vector(19 downto 0); -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_mem_address -> intel_generic_serial_flash_interface_top_0:avl_mem_address
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_read          : std_logic;                     -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_mem_read -> intel_generic_serial_flash_interface_top_0:avl_mem_read
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_mem_byteenable -> intel_generic_serial_flash_interface_top_0:avl_mem_byteenable
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid : std_logic;                     -- intel_generic_serial_flash_interface_top_0:avl_mem_readdatavalid -> mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_write         : std_logic;                     -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_mem_write -> intel_generic_serial_flash_interface_top_0:avl_mem_write
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_mem_writedata -> intel_generic_serial_flash_interface_top_0:avl_mem_writedata
	signal mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_burstcount    : std_logic_vector(6 downto 0);  -- mm_interconnect_0:intel_generic_serial_flash_interface_top_0_avl_mem_burstcount -> intel_generic_serial_flash_interface_top_0:avl_mem_burstcount
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata                              : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata                            : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest                         : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess                         : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address                             : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                                : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                               : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                                     : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                                      : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                                        : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                                        : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_angle_barre_s1_chipselect                                        : std_logic;                     -- mm_interconnect_0:angle_barre_s1_chipselect -> angle_barre:chipselect
	signal mm_interconnect_0_angle_barre_s1_readdata                                          : std_logic_vector(31 downto 0); -- angle_barre:readdata -> mm_interconnect_0:angle_barre_s1_readdata
	signal mm_interconnect_0_angle_barre_s1_address                                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:angle_barre_s1_address -> angle_barre:address
	signal mm_interconnect_0_angle_barre_s1_write                                             : std_logic;                     -- mm_interconnect_0:angle_barre_s1_write -> mm_interconnect_0_angle_barre_s1_write:in
	signal mm_interconnect_0_angle_barre_s1_writedata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:angle_barre_s1_writedata -> angle_barre:writedata
	signal mm_interconnect_0_write_n_s1_readdata                                              : std_logic_vector(31 downto 0); -- write_n:readdata -> mm_interconnect_0:write_n_s1_readdata
	signal mm_interconnect_0_write_n_s1_address                                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:write_n_s1_address -> write_n:address
	signal mm_interconnect_0_write_data_s1_readdata                                           : std_logic_vector(31 downto 0); -- write_data:readdata -> mm_interconnect_0:write_data_s1_readdata
	signal mm_interconnect_0_write_data_s1_address                                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:write_data_s1_address -> write_data:address
	signal mm_interconnect_0_butee_g_s1_chipselect                                            : std_logic;                     -- mm_interconnect_0:butee_g_s1_chipselect -> butee_g:chipselect
	signal mm_interconnect_0_butee_g_s1_readdata                                              : std_logic_vector(31 downto 0); -- butee_g:readdata -> mm_interconnect_0:butee_g_s1_readdata
	signal mm_interconnect_0_butee_g_s1_address                                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:butee_g_s1_address -> butee_g:address
	signal mm_interconnect_0_butee_g_s1_write                                                 : std_logic;                     -- mm_interconnect_0:butee_g_s1_write -> mm_interconnect_0_butee_g_s1_write:in
	signal mm_interconnect_0_butee_g_s1_writedata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:butee_g_s1_writedata -> butee_g:writedata
	signal mm_interconnect_0_butee_d_s1_chipselect                                            : std_logic;                     -- mm_interconnect_0:butee_d_s1_chipselect -> butee_d:chipselect
	signal mm_interconnect_0_butee_d_s1_readdata                                              : std_logic_vector(31 downto 0); -- butee_d:readdata -> mm_interconnect_0:butee_d_s1_readdata
	signal mm_interconnect_0_butee_d_s1_address                                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:butee_d_s1_address -> butee_d:address
	signal mm_interconnect_0_butee_d_s1_write                                                 : std_logic;                     -- mm_interconnect_0:butee_d_s1_write -> mm_interconnect_0_butee_d_s1_write:in
	signal mm_interconnect_0_butee_d_s1_writedata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:butee_d_s1_writedata -> butee_d:writedata
	signal mm_interconnect_0_freq_s1_chipselect                                               : std_logic;                     -- mm_interconnect_0:freq_s1_chipselect -> freq:chipselect
	signal mm_interconnect_0_freq_s1_readdata                                                 : std_logic_vector(31 downto 0); -- freq:readdata -> mm_interconnect_0:freq_s1_readdata
	signal mm_interconnect_0_freq_s1_address                                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:freq_s1_address -> freq:address
	signal mm_interconnect_0_freq_s1_write                                                    : std_logic;                     -- mm_interconnect_0:freq_s1_write -> mm_interconnect_0_freq_s1_write:in
	signal mm_interconnect_0_freq_s1_writedata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:freq_s1_writedata -> freq:writedata
	signal mm_interconnect_0_duty_s1_chipselect                                               : std_logic;                     -- mm_interconnect_0:duty_s1_chipselect -> duty:chipselect
	signal mm_interconnect_0_duty_s1_readdata                                                 : std_logic_vector(31 downto 0); -- duty:readdata -> mm_interconnect_0:duty_s1_readdata
	signal mm_interconnect_0_duty_s1_address                                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:duty_s1_address -> duty:address
	signal mm_interconnect_0_duty_s1_write                                                    : std_logic;                     -- mm_interconnect_0:duty_s1_write -> mm_interconnect_0_duty_s1_write:in
	signal mm_interconnect_0_duty_s1_writedata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:duty_s1_writedata -> duty:writedata
	signal mm_interconnect_0_sens_s1_chipselect                                               : std_logic;                     -- mm_interconnect_0:sens_s1_chipselect -> sens:chipselect
	signal mm_interconnect_0_sens_s1_readdata                                                 : std_logic_vector(31 downto 0); -- sens:readdata -> mm_interconnect_0:sens_s1_readdata
	signal mm_interconnect_0_sens_s1_address                                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sens_s1_address -> sens:address
	signal mm_interconnect_0_sens_s1_write                                                    : std_logic;                     -- mm_interconnect_0:sens_s1_write -> mm_interconnect_0_sens_s1_write:in
	signal mm_interconnect_0_sens_s1_writedata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:sens_s1_writedata -> sens:writedata
	signal irq_mapper_receiver0_irq                                                           : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal nios2_gen2_0_irq_irq                                                               : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                                     : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:intel_generic_serial_flash_interface_top_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                                 : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                                 : std_logic;                     -- rst_controller_001:reset_out -> intel_generic_serial_flash_interface_top_0:reset_reset
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv                     : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_angle_barre_s1_write_ports_inv                                   : std_logic;                     -- mm_interconnect_0_angle_barre_s1_write:inv -> angle_barre:write_n
	signal mm_interconnect_0_butee_g_s1_write_ports_inv                                       : std_logic;                     -- mm_interconnect_0_butee_g_s1_write:inv -> butee_g:write_n
	signal mm_interconnect_0_butee_d_s1_write_ports_inv                                       : std_logic;                     -- mm_interconnect_0_butee_d_s1_write:inv -> butee_d:write_n
	signal mm_interconnect_0_freq_s1_write_ports_inv                                          : std_logic;                     -- mm_interconnect_0_freq_s1_write:inv -> freq:write_n
	signal mm_interconnect_0_duty_s1_write_ports_inv                                          : std_logic;                     -- mm_interconnect_0_duty_s1_write:inv -> duty:write_n
	signal mm_interconnect_0_sens_s1_write_ports_inv                                          : std_logic;                     -- mm_interconnect_0_sens_s1_write:inv -> sens:write_n
	signal rst_controller_reset_out_reset_ports_inv                                           : std_logic;                     -- rst_controller_reset_out_reset:inv -> [angle_barre:reset_n, butee_d:reset_n, butee_g:reset_n, duty:reset_n, freq:reset_n, jtag_uart_0:rst_n, nios2_gen2_0:reset_n, sens:reset_n, sysid_qsys_0:reset_n, write_data:reset_n, write_n:reset_n]

begin

	angle_barre : component sopc3_angle_barre
		port map (
			clk        => clk_clk,                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_angle_barre_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_angle_barre_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_angle_barre_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_angle_barre_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_angle_barre_s1_readdata,        --                    .readdata
			out_port   => angle_barre_external_connection_export            -- external_connection.export
		);

	butee_d : component sopc3_angle_barre
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_butee_d_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_butee_d_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_butee_d_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_butee_d_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_butee_d_s1_readdata,        --                    .readdata
			out_port   => butee_d_external_connection_export            -- external_connection.export
		);

	butee_g : component sopc3_angle_barre
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_butee_g_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_butee_g_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_butee_g_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_butee_g_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_butee_g_s1_readdata,        --                    .readdata
			out_port   => butee_g_external_connection_export            -- external_connection.export
		);

	duty : component sopc3_duty
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_duty_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_duty_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_duty_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_duty_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_duty_s1_readdata,        --                    .readdata
			out_port   => duty_external_connection_export            -- external_connection.export
		);

	freq : component sopc3_duty
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_freq_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_freq_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_freq_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_freq_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_freq_s1_readdata,        --                    .readdata
			out_port   => freq_external_connection_export            -- external_connection.export
		);

	intel_generic_serial_flash_interface_top_0 : component sopc3_intel_generic_serial_flash_interface_top_0
		generic map (
			DEVICE_FAMILY => "Cyclone IV E",
			CHIP_SELS     => 1
		)
		port map (
			avl_csr_address       => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_address,       -- avl_csr.address
			avl_csr_read          => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_read,          --        .read
			avl_csr_readdata      => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_readdata,      --        .readdata
			avl_csr_write         => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_write,         --        .write
			avl_csr_writedata     => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_writedata,     --        .writedata
			avl_csr_waitrequest   => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest,   --        .waitrequest
			avl_csr_readdatavalid => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid, --        .readdatavalid
			avl_mem_write         => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_write,         -- avl_mem.write
			avl_mem_burstcount    => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_burstcount,    --        .burstcount
			avl_mem_waitrequest   => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest,   --        .waitrequest
			avl_mem_read          => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_read,          --        .read
			avl_mem_address       => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_address,       --        .address
			avl_mem_writedata     => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_writedata,     --        .writedata
			avl_mem_readdata      => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_readdata,      --        .readdata
			avl_mem_readdatavalid => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid, --        .readdatavalid
			avl_mem_byteenable    => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_byteenable,    --        .byteenable
			clk_clk               => clk_clk,                                                                            --     clk.clk
			reset_reset           => rst_controller_001_reset_out_reset                                                  --   reset.reset
		);

	jtag_uart_0 : component sopc3_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	nios2_gen2_0 : component sopc3_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component sopc3_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	sens : component sopc3_sens
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_sens_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_sens_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_sens_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_sens_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_sens_s1_readdata,        --                    .readdata
			out_port   => sens_external_connection_export            -- external_connection.export
		);

	sysid_qsys_0 : component sopc3_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	write_data : component sopc3_write_data
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_write_data_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_write_data_s1_readdata, --                    .readdata
			in_port  => write_data_external_connection_export     -- external_connection.export
		);

	write_n : component sopc3_write_n
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_write_n_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_write_n_s1_readdata,    --                    .readdata
			in_port  => write_n_external_connection_export        -- external_connection.export
		);

	mm_interconnect_0 : component sopc3_mm_interconnect_0
		port map (
			clk_0_clk_clk                                                                => clk_clk,                                                                            --                                                              clk_0_clk.clk
			intel_generic_serial_flash_interface_top_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                                     -- intel_generic_serial_flash_interface_top_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                               => rst_controller_reset_out_reset,                                                     --                               nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                                             => nios2_gen2_0_data_master_address,                                                   --                                               nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                                         => nios2_gen2_0_data_master_waitrequest,                                               --                                                                       .waitrequest
			nios2_gen2_0_data_master_byteenable                                          => nios2_gen2_0_data_master_byteenable,                                                --                                                                       .byteenable
			nios2_gen2_0_data_master_read                                                => nios2_gen2_0_data_master_read,                                                      --                                                                       .read
			nios2_gen2_0_data_master_readdata                                            => nios2_gen2_0_data_master_readdata,                                                  --                                                                       .readdata
			nios2_gen2_0_data_master_write                                               => nios2_gen2_0_data_master_write,                                                     --                                                                       .write
			nios2_gen2_0_data_master_writedata                                           => nios2_gen2_0_data_master_writedata,                                                 --                                                                       .writedata
			nios2_gen2_0_data_master_debugaccess                                         => nios2_gen2_0_data_master_debugaccess,                                               --                                                                       .debugaccess
			nios2_gen2_0_instruction_master_address                                      => nios2_gen2_0_instruction_master_address,                                            --                                        nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                                  => nios2_gen2_0_instruction_master_waitrequest,                                        --                                                                       .waitrequest
			nios2_gen2_0_instruction_master_read                                         => nios2_gen2_0_instruction_master_read,                                               --                                                                       .read
			nios2_gen2_0_instruction_master_readdata                                     => nios2_gen2_0_instruction_master_readdata,                                           --                                                                       .readdata
			angle_barre_s1_address                                                       => mm_interconnect_0_angle_barre_s1_address,                                           --                                                         angle_barre_s1.address
			angle_barre_s1_write                                                         => mm_interconnect_0_angle_barre_s1_write,                                             --                                                                       .write
			angle_barre_s1_readdata                                                      => mm_interconnect_0_angle_barre_s1_readdata,                                          --                                                                       .readdata
			angle_barre_s1_writedata                                                     => mm_interconnect_0_angle_barre_s1_writedata,                                         --                                                                       .writedata
			angle_barre_s1_chipselect                                                    => mm_interconnect_0_angle_barre_s1_chipselect,                                        --                                                                       .chipselect
			butee_d_s1_address                                                           => mm_interconnect_0_butee_d_s1_address,                                               --                                                             butee_d_s1.address
			butee_d_s1_write                                                             => mm_interconnect_0_butee_d_s1_write,                                                 --                                                                       .write
			butee_d_s1_readdata                                                          => mm_interconnect_0_butee_d_s1_readdata,                                              --                                                                       .readdata
			butee_d_s1_writedata                                                         => mm_interconnect_0_butee_d_s1_writedata,                                             --                                                                       .writedata
			butee_d_s1_chipselect                                                        => mm_interconnect_0_butee_d_s1_chipselect,                                            --                                                                       .chipselect
			butee_g_s1_address                                                           => mm_interconnect_0_butee_g_s1_address,                                               --                                                             butee_g_s1.address
			butee_g_s1_write                                                             => mm_interconnect_0_butee_g_s1_write,                                                 --                                                                       .write
			butee_g_s1_readdata                                                          => mm_interconnect_0_butee_g_s1_readdata,                                              --                                                                       .readdata
			butee_g_s1_writedata                                                         => mm_interconnect_0_butee_g_s1_writedata,                                             --                                                                       .writedata
			butee_g_s1_chipselect                                                        => mm_interconnect_0_butee_g_s1_chipselect,                                            --                                                                       .chipselect
			duty_s1_address                                                              => mm_interconnect_0_duty_s1_address,                                                  --                                                                duty_s1.address
			duty_s1_write                                                                => mm_interconnect_0_duty_s1_write,                                                    --                                                                       .write
			duty_s1_readdata                                                             => mm_interconnect_0_duty_s1_readdata,                                                 --                                                                       .readdata
			duty_s1_writedata                                                            => mm_interconnect_0_duty_s1_writedata,                                                --                                                                       .writedata
			duty_s1_chipselect                                                           => mm_interconnect_0_duty_s1_chipselect,                                               --                                                                       .chipselect
			freq_s1_address                                                              => mm_interconnect_0_freq_s1_address,                                                  --                                                                freq_s1.address
			freq_s1_write                                                                => mm_interconnect_0_freq_s1_write,                                                    --                                                                       .write
			freq_s1_readdata                                                             => mm_interconnect_0_freq_s1_readdata,                                                 --                                                                       .readdata
			freq_s1_writedata                                                            => mm_interconnect_0_freq_s1_writedata,                                                --                                                                       .writedata
			freq_s1_chipselect                                                           => mm_interconnect_0_freq_s1_chipselect,                                               --                                                                       .chipselect
			intel_generic_serial_flash_interface_top_0_avl_csr_address                   => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_address,       --                     intel_generic_serial_flash_interface_top_0_avl_csr.address
			intel_generic_serial_flash_interface_top_0_avl_csr_write                     => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_write,         --                                                                       .write
			intel_generic_serial_flash_interface_top_0_avl_csr_read                      => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_read,          --                                                                       .read
			intel_generic_serial_flash_interface_top_0_avl_csr_readdata                  => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_readdata,      --                                                                       .readdata
			intel_generic_serial_flash_interface_top_0_avl_csr_writedata                 => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_writedata,     --                                                                       .writedata
			intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid             => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_readdatavalid, --                                                                       .readdatavalid
			intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest               => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_csr_waitrequest,   --                                                                       .waitrequest
			intel_generic_serial_flash_interface_top_0_avl_mem_address                   => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_address,       --                     intel_generic_serial_flash_interface_top_0_avl_mem.address
			intel_generic_serial_flash_interface_top_0_avl_mem_write                     => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_write,         --                                                                       .write
			intel_generic_serial_flash_interface_top_0_avl_mem_read                      => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_read,          --                                                                       .read
			intel_generic_serial_flash_interface_top_0_avl_mem_readdata                  => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_readdata,      --                                                                       .readdata
			intel_generic_serial_flash_interface_top_0_avl_mem_writedata                 => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_writedata,     --                                                                       .writedata
			intel_generic_serial_flash_interface_top_0_avl_mem_burstcount                => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_burstcount,    --                                                                       .burstcount
			intel_generic_serial_flash_interface_top_0_avl_mem_byteenable                => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_byteenable,    --                                                                       .byteenable
			intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid             => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_readdatavalid, --                                                                       .readdatavalid
			intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest               => mm_interconnect_0_intel_generic_serial_flash_interface_top_0_avl_mem_waitrequest,   --                                                                       .waitrequest
			jtag_uart_0_avalon_jtag_slave_address                                        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,                            --                                          jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                                          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                              --                                                                       .write
			jtag_uart_0_avalon_jtag_slave_read                                           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                               --                                                                       .read
			jtag_uart_0_avalon_jtag_slave_readdata                                       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,                           --                                                                       .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                                      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,                          --                                                                       .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,                        --                                                                       .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,                         --                                                                       .chipselect
			nios2_gen2_0_debug_mem_slave_address                                         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,                             --                                           nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                                           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                               --                                                                       .write
			nios2_gen2_0_debug_mem_slave_read                                            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                                --                                                                       .read
			nios2_gen2_0_debug_mem_slave_readdata                                        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,                            --                                                                       .readdata
			nios2_gen2_0_debug_mem_slave_writedata                                       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,                           --                                                                       .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                                      => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,                          --                                                                       .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,                         --                                                                       .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,                         --                                                                       .debugaccess
			onchip_memory2_0_s1_address                                                  => mm_interconnect_0_onchip_memory2_0_s1_address,                                      --                                                    onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                                    => mm_interconnect_0_onchip_memory2_0_s1_write,                                        --                                                                       .write
			onchip_memory2_0_s1_readdata                                                 => mm_interconnect_0_onchip_memory2_0_s1_readdata,                                     --                                                                       .readdata
			onchip_memory2_0_s1_writedata                                                => mm_interconnect_0_onchip_memory2_0_s1_writedata,                                    --                                                                       .writedata
			onchip_memory2_0_s1_byteenable                                               => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                                   --                                                                       .byteenable
			onchip_memory2_0_s1_chipselect                                               => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                                   --                                                                       .chipselect
			onchip_memory2_0_s1_clken                                                    => mm_interconnect_0_onchip_memory2_0_s1_clken,                                        --                                                                       .clken
			sens_s1_address                                                              => mm_interconnect_0_sens_s1_address,                                                  --                                                                sens_s1.address
			sens_s1_write                                                                => mm_interconnect_0_sens_s1_write,                                                    --                                                                       .write
			sens_s1_readdata                                                             => mm_interconnect_0_sens_s1_readdata,                                                 --                                                                       .readdata
			sens_s1_writedata                                                            => mm_interconnect_0_sens_s1_writedata,                                                --                                                                       .writedata
			sens_s1_chipselect                                                           => mm_interconnect_0_sens_s1_chipselect,                                               --                                                                       .chipselect
			sysid_qsys_0_control_slave_address                                           => mm_interconnect_0_sysid_qsys_0_control_slave_address,                               --                                             sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                                          => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,                              --                                                                       .readdata
			write_data_s1_address                                                        => mm_interconnect_0_write_data_s1_address,                                            --                                                          write_data_s1.address
			write_data_s1_readdata                                                       => mm_interconnect_0_write_data_s1_readdata,                                           --                                                                       .readdata
			write_n_s1_address                                                           => mm_interconnect_0_write_n_s1_address,                                               --                                                             write_n_s1.address
			write_n_s1_readdata                                                          => mm_interconnect_0_write_n_s1_readdata                                               --                                                                       .readdata
		);

	irq_mapper : component sopc3_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component sopc3_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component sopc3_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => open,                                   --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_angle_barre_s1_write_ports_inv <= not mm_interconnect_0_angle_barre_s1_write;

	mm_interconnect_0_butee_g_s1_write_ports_inv <= not mm_interconnect_0_butee_g_s1_write;

	mm_interconnect_0_butee_d_s1_write_ports_inv <= not mm_interconnect_0_butee_d_s1_write;

	mm_interconnect_0_freq_s1_write_ports_inv <= not mm_interconnect_0_freq_s1_write;

	mm_interconnect_0_duty_s1_write_ports_inv <= not mm_interconnect_0_duty_s1_write;

	mm_interconnect_0_sens_s1_write_ports_inv <= not mm_interconnect_0_sens_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of sopc3
